parameter N = 4;