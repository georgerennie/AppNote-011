`define IDX0 2